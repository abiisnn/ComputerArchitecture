LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ROM IS
	-- VALORES GENERICOS DE LA MEMORIA DE PROGRAMA DEL ESCOMIPS
	GENERIC (
		BITS_D : INTEGER := 25;
		BITS_A : INTEGER := 16);

	-- PUERTOS DE ENTRADA (BUS DE DIRECCIONES 'A')
	-- Y SALIDA (BUS DE DIRECCIONES 'D')
    PORT (
		A : IN STD_LOGIC_VECTOR (BITS_A - 1 DOWNTO 0);
		D : OUT STD_LOGIC_VECTOR (BITS_D - 1 DOWNTO 0));
END ROM;

ARCHITECTURE FUNCIONAMIENTO OF ROM IS
	
	-- DEFINICI�N DEL TIPO DE DATO MEMORIA
	TYPE MEMORIA IS ARRAY (0 TO 2 ** BITS_A - 1) 
		OF STD_LOGIC_VECTOR(BITS_D - 1 DOWNTO 0); 

	-- DECLARACI�N DE UNA MEMORIA ROM CON EL PROGRAMA DE EJEMPLO.
	CONSTANT ROM : MEMORIA := (
		"0000100000000000000010111",
		"0001100000000000000001010",
		"0000100000000000010000010",
		"0001100000000000000001011",
		"0000100000000000001000110",
		"0001100000000000000001100",
		"0000100000000000100000100",
		"0001100000000000000001101",
		"0000100001111111111010011",
		"0001100000000000000001110",
		"0000100000000000010110100",
		"0001100000000000000001111",
		"0000100000000000000000000",
		"0000100010000000000000000",
		"0000100100000000000000000",
		"0000100110000000000000110",
		"0011001000011000000000001",
		"1001001000000000000001110",
		"0000100010000000000000000",
		"0000001010100000000000001",
		"1001001010001000000001001",
		"1011101100001000000001010",
		"1011101110001000000001011",
		"1000001110110000000000100",
		"1011100100001000000001010",
		"0010001110001000000001010",
		"0010000100001000000001011",
		"0010100010001000000000001",
		"1001100000000000000010100",
		"0010100000000000000000001",
		"1001100000000000000010001",
		"1011000000000000000000000",
		"1001100000000000000011111",
		OTHERS => (OTHERS => '0'));

BEGIN

	D <= ROM(CONV_INTEGER(A));


END FUNCIONAMIENTO;

