	
	stim_proc: process
	begin
		DATAIN <= "10010101";
		SHIFT <= "100"
	wait for 100 ns;

		wait;
	end process;