library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity mem_funcion is
    Port ( FUNCODE : in  STD_LOGIC_VECTOR (3 downto 0);
           MICROINSTRUCCION : out  STD_LOGIC_VECTOR (19 downto 0));
end mem_funcion;

architecture Behavioral of mem_funcion is

type memoria is array (0 to 15) of std_logic_vector(19 downto 0);
constant rom: memoria := (
	"00000100110000011001", --00 ADD
	"00000100110000111001", --01 SUB
	"00000100110000000001", --02 AND
	"00000100110000001001", --03 OR
	"00000100110000010001", --04 XOR
	"00000100110001101001", --05 NAND
	"00000100110001100001", --06 NOR
	"00000100110001010001", --07 XNOR
	"00000100110001101001", --08 NOT
	"00000011000000000000", --09 SLL
	"00000010000000000000", --10 SRL
	"00000000000000000000", --11
	"00000000000000000000", --12
	"00000000000000000000", --13
	"00000000000000000000", --14
	"00000000000000000000"  --15
);

begin

	MICROINSTRUCCION <= rom(conv_integer(FUNCODE));

end Behavioral;

