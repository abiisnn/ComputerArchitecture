library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity mem_operacion is
    Port ( OPCODE : in  STD_LOGIC_VECTOR (4 downto 0);
           MICROINSTRUCCION : out  STD_LOGIC_VECTOR (19 downto 0));
end mem_operacion;

architecture Behavioral of mem_operacion is

type memoria is array (0 to 31) of std_logic_vector(19 downto 0);
constant rom: memoria := (
	"00001000010000111000", --00 Bcond
	"00000000100000000000", --01 LI
	"00000100100000000100", --02 LWI
	"00001000000000000110", --03 SWI
	"00001000001010011010", --04 SW
	"00000100110010011001", --05 ADDI
	"00000100110010111001", --06 SUBI
	"00000100111010000001", --07 ANDI
	"00000100111010001001", --08 ORI
	"00000100111010010001", --09 XORI
	"00000100111011101001", --10 NANDI
	"00000100111011100001", --11 NORI
	"00000100111011010001", --12 XNORI
	"00110000000110011001", --13 BEQI
	"00110000000110011001", --14 BNEI
	"00110000000110011001", --15 BLTI
	"00110000000110011001", --16 BLETI
	"00110000000110011001", --17 BGTI
	"00110000000110011001", --18 BGETI
	"00100000000000000000", --19 B
	"10100000000000000000", --20 CALL
	"01100000000000000000", --21 RET
	"00000000000000000000", --22 NOP
	"00000100101010011000", --23 LW
	"00000000000000000000", --24
	"00000000000000000000", --25
	"00000000000000000000", --26
	"00000000000000000000", --27
	"00000000000000000000", --28
	"00000000000000000000", --29
	"00000000000000000000", --30
	"00000000000000000000"  --31
);

begin

	MICROINSTRUCCION <= rom(conv_integer(OPCODE));

end Behavioral;

